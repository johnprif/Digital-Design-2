library ieee;
use ieee.std_logic_1164.all;

package Declarations is
		type state_type is (LOAD, ADD, SHIFT, FINISH);
end Declarations;

